package fifo_package;
    `include "fifo_transaction.sv"
    `include "fifo_generator.sv"
    `include "fifo_driver.sv"
    `include "fifo_enviroment.sv"
    `include "fifo_test.sv"
endpackage